module and_logic(
  input A, B,
  output Y
);

  assign Y = A & B;

endmodule
  
