module or_logic(
  input A, B,
  output Y
);

  assign Y = A | B;

endmodule
  
